`define CLW32
//`define MR
//`define TWO

